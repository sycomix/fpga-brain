altfpcompM_inst : altfpcompM PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		agb	 => agb_sig
	);
