altfpcomp_inst : altfpcomp PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		alb	 => alb_sig
	);
