library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
ENTITY VGA IS
PORT(
	CLOCK_INVGA: IN STD_LOGIC;
	netOuts: IN STD_LOGIC_VECTOR(15 downto 0);
	VGA_HS, VGA_VS: OUT STD_LOGIC;
	VGA_R, VGA_G, VGA_B: OUT STD_LOGIC;
	vgaTick: OUT STD_LOGIC
);
END VGA;
 
ARCHITECTURE MAIN OF VGA IS
 
COMPONENT SYNC IS
PORT(
	CLK: IN STD_LOGIC;
	netOuts: IN STD_LOGIC_VECTOR(15 downto 0);
	HSYNC, VSYNC: OUT STD_LOGIC;
	R, G, B: OUT STD_LOGIC;
	vgaTick: OUT STD_LOGIC
);
END COMPONENT SYNC;
 
BEGIN
C1: SYNC PORT MAP (CLOCK_INVGA, netOuts, VGA_HS, VGA_VS, VGA_R, VGA_G, VGA_B, vgaTick);
 
END ARCHITECTURE MAIN;
